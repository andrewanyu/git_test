class vseq extends uvm_sequence;

this this this 

haha;

super super super

function new();
    hahah;
    
endfunction


endclass: vseq
