class vseq extends uvm_sequence;

this this this 

super super super

  function new();
  endfunction: new

endclass: vseq
