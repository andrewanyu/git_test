class vseq extends uvm_sequence;

this this this 

super super super



endclass: vseq